
module clk_div2(input clk, input reset, output reg clk_out);
    always @(posedge clk or posedge reset) begin
        if (reset) clk_out <= 1'b0;
        else       clk_out <= ~clk_out;
    end
endmodule
